`timescale 1ps/1ps

module Pipe_Line_Test_Bench ();
    
endmodule