module IF_Stage (
    input clk, rst, freeze, Branch_taken,
    input [31:0]BranchAddr,
    output [31:0]PC, Instruction
);
    
endmodule