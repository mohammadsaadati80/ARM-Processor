module Pipe_Line_Test_Bench ();
    
endmodule