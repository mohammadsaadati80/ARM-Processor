module Instruction_mem (
    input clk, rst,
    input [31:0]PC,
    output reg [31:0]Instruction
);

    // ¯\_(ツ)_/¯
    
endmodule